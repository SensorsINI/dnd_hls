// This file is part of https://github.com/SensorsINI/dnd_hls. 
// This intellectual property is licensed under the terms of the project license available at the root of the project.

`timescale 1ns/1ps

module luts #(N1=98, N2=10)(
  output wire [N2-1:0][N1/2:0][6-1:0] weights_n1_mag,
  output wire [N2-1:0][N1/2:0][6-1:0] weights_n1_pol,
  output wire [N2  :0][4-1:0] weights_n2
);
  assign weights_n1_mag = '{
    '{  6'd8     ,  6'd0     , -6'd6     ,  6'd6     , -6'd4     ,  6'd0     ,  6'd0     ,  6'd0     ,  6'd2     ,  6'd4     ,  6'd10    ,  6'd0     ,  6'd2     ,  6'd4     ,  6'd6     ,  6'd4     ,  6'd6     ,  6'd2     ,  6'd0     ,  6'd12    ,  6'd0     ,  6'd0     ,  6'd2     , -6'd4     ,  6'd0     , -6'd14    ,  6'd0     , -6'd2     , -6'd2     ,  6'd0     ,  6'd0     ,  6'd10    ,  6'd2     ,  6'd10    ,  6'd6     ,  6'd0     ,  6'd0     ,  6'd0     ,  6'd10    , -6'd4     ,  6'd2     ,  6'd2     ,  6'd6     ,  6'd6     , -6'd4     ,  6'd0     , -6'd4     ,  6'd4     , -6'd2     ,  6'd6      },
    '{ -6'd8     , -6'd2     ,  6'd4     ,  6'd4     , -6'd2     ,  6'd2     , -6'd8     , -6'd6     ,  6'd0     , -6'd4     ,  6'd4     ,  6'd0     ,  6'd0     ,  6'd0     ,  6'd4     , -6'd2     ,  6'd6     , -6'd6     ,  6'd0     , -6'd6     ,  6'd2     ,  6'd6     ,  6'd0     ,  6'd2     , -6'd8     ,  6'd0     , -6'd8     ,  6'd6     , -6'd6     ,  6'd2     ,  6'd0     ,  6'd4     , -6'd14    , -6'd2     , -6'd4     ,  6'd8     , -6'd8     ,  6'd6     ,  6'd2     ,  6'd10    ,  6'd2     ,  6'd2     , -6'd2     , -6'd6     , -6'd2     , -6'd4     , -6'd6     , -6'd2     , -6'd4     , -6'd6      },
    '{  6'd8     ,  6'd10    ,  6'd10    , -6'd4     , -6'd8     , -6'd8     , -6'd4     ,  6'd4     ,  6'd2     ,  6'd6     , -6'd6     , -6'd10    , -6'd2     , -6'd2     , -6'd4     , -6'd2     ,  6'd4     ,  6'd0     , -6'd14    , -6'd4     , -6'd2     ,  6'd2     , -6'd6     ,  6'd4     , -6'd4     , -6'd6     , -6'd6     ,  6'd0     , -6'd6     , -6'd4     , -6'd4     ,  6'd0     , -6'd8     , -6'd2     , -6'd4     , -6'd2     , -6'd6     ,  6'd0     , -6'd4     , -6'd10    , -6'd8     ,  6'd0     , -6'd4     , -6'd8     ,  6'd2     ,  6'd2     , -6'd10    , -6'd4     , -6'd6     , -6'd6      },
    '{ -6'd16    ,  6'd0     ,  6'd4     ,  6'd4     ,  6'd0     ,  6'd1     , -6'd2     , -6'd3     ,  6'd0     , -6'd2     ,  6'd5     ,  6'd0     ,  6'd7     ,  6'd5     ,  6'd3     ,  6'd3     ,  6'd2     ,  6'd3     ,  6'd6     ,  6'd3     ,  6'd2     ,  6'd4     ,  6'd2     ,  6'd3     ,  6'd6     , -6'd3     ,  6'd3     ,  6'd0     ,  6'd1     ,  6'd2     ,  6'd1     ,  6'd6     ,  6'd6     ,  6'd1     ,  6'd2     , -6'd1     , -6'd2     ,  6'd2     ,  6'd1     ,  6'd3     ,  6'd2     ,  6'd1     , -6'd6     , -6'd1     ,  6'd3     ,  6'd3     ,  6'd4     , -6'd3     ,  6'd1     , -6'd1      },
    '{ -6'd8     , -6'd2     , -6'd4     ,  6'd2     , -6'd2     ,  6'd2     , -6'd2     ,  6'd0     , -6'd2     , -6'd6     ,  6'd2     ,  6'd2     , -6'd2     , -6'd6     , -6'd2     ,  6'd2     ,  6'd0     ,  6'd0     , -6'd2     , -6'd8     ,  6'd2     , -6'd2     , -6'd4     , -6'd2     ,  6'd2     ,  6'd6     ,  6'd6     , -6'd8     , -6'd6     ,  6'd4     , -6'd6     , -6'd4     , -6'd8     , -6'd2     , -6'd2     , -6'd4     ,  6'd6     , -6'd4     ,  6'd0     ,  6'd4     , -6'd6     ,  6'd4     ,  6'd0     , -6'd2     , -6'd6     ,  6'd2     , -6'd6     , -6'd6     ,  6'd4     , -6'd4      },
    '{  6'd8     , -6'd2     , -6'd4     , -6'd2     ,  6'd0     , -6'd4     , -6'd2     , -6'd2     ,  6'd0     ,  6'd2     ,  6'd2     ,  6'd0     ,  6'd6     ,  6'd0     ,  6'd10    ,  6'd0     , -6'd4     ,  6'd0     ,  6'd6     ,  6'd0     ,  6'd8     ,  6'd8     , -6'd4     ,  6'd0     ,  6'd6     , -6'd8     , -6'd4     , -6'd4     ,  6'd4     ,  6'd4     ,  6'd0     ,  6'd6     ,  6'd10    ,  6'd2     , -6'd12    ,  6'd0     ,  6'd8     , -6'd8     ,  6'd2     ,  6'd8     , -6'd4     , -6'd10    ,  6'd2     ,  6'd0     ,  6'd6     , -6'd4     ,  6'd6     ,  6'd0     , -6'd8     ,  6'd8      },
    '{  6'd0     ,  6'd2     , -6'd4     ,  6'd0     ,  6'd2     ,  6'd8     ,  6'd0     , -6'd4     ,  6'd8     , -6'd2     , -6'd2     ,  6'd0     , -6'd2     , -6'd4     , -6'd2     ,  6'd2     , -6'd4     ,  6'd0     ,  6'd12    ,  6'd2     , -6'd2     ,  6'd2     , -6'd2     ,  6'd6     ,  6'd8     , -6'd4     ,  6'd6     ,  6'd6     , -6'd2     ,  6'd2     ,  6'd0     ,  6'd2     ,  6'd4     ,  6'd6     ,  6'd2     ,  6'd0     ,  6'd4     ,  6'd4     , -6'd4     ,  6'd0     ,  6'd6     ,  6'd0     ,  6'd0     , -6'd2     ,  6'd2     ,  6'd2     ,  6'd4     , -6'd2     ,  6'd4     , -6'd4      },
    '{  6'd0     , -6'd6     ,  6'd0     ,  6'd8     ,  6'd4     , -6'd4     ,  6'd4     ,  6'd0     , -6'd6     ,  6'd6     ,  6'd0     ,  6'd8     , -6'd2     , -6'd2     ,  6'd2     , -6'd4     ,  6'd0     ,  6'd2     ,  6'd2     , -6'd2     , -6'd4     ,  6'd6     ,  6'd6     ,  6'd6     ,  6'd6     , -6'd14    ,  6'd4     ,  6'd8     ,  6'd4     ,  6'd2     ,  6'd8     ,  6'd0     ,  6'd4     ,  6'd8     , -6'd4     ,  6'd2     , -6'd6     , -6'd4     , -6'd2     ,  6'd10    ,  6'd4     ,  6'd6     , -6'd2     , -6'd6     , -6'd6     ,  6'd2     ,  6'd6     , -6'd2     , -6'd4     , -6'd2      },
    '{  6'd0     , -6'd2     , -6'd2     ,  6'd2     ,  6'd0     , -6'd2     , -6'd4     , -6'd2     ,  6'd0     ,  6'd0     ,  6'd2     , -6'd8     ,  6'd4     ,  6'd2     , -6'd2     ,  6'd0     ,  6'd0     , -6'd2     ,  6'd0     , -6'd4     ,  6'd4     ,  6'd2     , -6'd4     ,  6'd2     ,  6'd2     ,  6'd0     , -6'd6     , -6'd2     , -6'd2     ,  6'd0     , -6'd4     ,  6'd0     ,  6'd0     ,  6'd4     , -6'd4     ,  6'd0     , -6'd4     ,  6'd0     , -6'd10    , -6'd8     , -6'd2     , -6'd2     , -6'd6     , -6'd2     , -6'd2     ,  6'd2     ,  6'd2     , -6'd4     ,  6'd0     ,  6'd4      },
    '{  6'd0     , -6'd6     , -6'd2     , -6'd6     , -6'd8     ,  6'd0     , -6'd2     ,  6'd4     , -6'd10    , -6'd2     , -6'd8     , -6'd10    ,  6'd0     , -6'd2     ,  6'd4     ,  6'd0     , -6'd2     ,  6'd2     , -6'd4     , -6'd6     ,  6'd10    ,  6'd6     , -6'd2     ,  6'd0     ,  6'd2     , -6'd6     ,  6'd4     ,  6'd8     ,  6'd2     ,  6'd2     ,  6'd0     , -6'd2     , -6'd4     , -6'd6     ,  6'd4     ,  6'd8     ,  6'd4     ,  6'd8     , -6'd6     , -6'd4     ,  6'd2     , -6'd2     , -6'd2     ,  6'd4     , -6'd6     , -6'd2     , -6'd4     , -6'd2     ,  6'd8     , -6'd2      }
  };

  assign weights_n1_pol = '{
    '{  6'd0     ,  6'd8     ,  6'd0     ,  6'd4     , -6'd2     ,  6'd2     ,  6'd2     ,  6'd2     , -6'd2     ,  6'd12    ,  6'd0     ,  6'd0     ,  6'd0     ,  6'd2     ,  6'd0     ,  6'd0     ,  6'd0     ,  6'd2     , -6'd2     ,  6'd4     ,  6'd2     ,  6'd4     , -6'd4     ,  6'd2     ,  6'd4     , -6'd14    ,  6'd2     ,  6'd4     , -6'd4     ,  6'd0     ,  6'd0     ,  6'd14    ,  6'd4     ,  6'd2     ,  6'd0     ,  6'd0     ,  6'd6     ,  6'd4     , -6'd6     , -6'd8     ,  6'd6     ,  6'd0     ,  6'd8     , -6'd4     ,  6'd2     ,  6'd2     ,  6'd0     ,  6'd6     ,  6'd0     , -6'd2      },
    '{  6'd0     , -6'd6     ,  6'd0     , -6'd2     , -6'd4     , -6'd2     ,  6'd0     ,  6'd0     ,  6'd0     ,  6'd2     ,  6'd0     , -6'd2     ,  6'd2     ,  6'd2     , -6'd6     , -6'd2     , -6'd2     , -6'd4     , -6'd4     , -6'd6     ,  6'd0     ,  6'd4     ,  6'd0     , -6'd6     , -6'd2     ,  6'd12    , -6'd8     ,  6'd6     , -6'd6     ,  6'd6     ,  6'd8     , -6'd2     , -6'd6     , -6'd2     , -6'd8     ,  6'd2     , -6'd4     , -6'd2     ,  6'd0     ,  6'd0     , -6'd4     ,  6'd6     ,  6'd2     , -6'd4     , -6'd4     , -6'd2     , -6'd4     ,  6'd0     , -6'd4     ,  6'd0      },
    '{  6'd0     ,  6'd0     , -6'd4     , -6'd4     ,  6'd10    ,  6'd0     ,  6'd0     ,  6'd0     , -6'd6     , -6'd2     ,  6'd4     ,  6'd8     ,  6'd4     , -6'd8     ,  6'd0     , -6'd4     ,  6'd0     , -6'd2     ,  6'd0     , -6'd6     , -6'd4     , -6'd2     ,  6'd2     , -6'd8     , -6'd2     , -6'd8     , -6'd8     , -6'd8     , -6'd8     , -6'd6     , -6'd4     , -6'd8     ,  6'd2     , -6'd4     ,  6'd2     ,  6'd4     , -6'd6     , -6'd4     ,  6'd2     ,  6'd6     ,  6'd0     ,  6'd10    ,  6'd4     ,  6'd0     ,  6'd0     ,  6'd2     ,  6'd4     , -6'd2     ,  6'd0     ,  6'd2      },
    '{  6'd0     ,  6'd2     , -6'd2     ,  6'd0     ,  6'd3     ,  6'd1     ,  6'd5     ,  6'd2     ,  6'd1     , -6'd2     ,  6'd3     ,  6'd2     ,  6'd0     ,  6'd2     ,  6'd3     ,  6'd3     ,  6'd1     , -6'd1     ,  6'd0     , -6'd1     ,  6'd0     ,  6'd0     ,  6'd0     , -6'd2     , -6'd1     ,  6'd1     , -6'd2     ,  6'd0     , -6'd4     , -6'd2     ,  6'd5     ,  6'd3     ,  6'd1     , -6'd2     ,  6'd1     ,  6'd2     ,  6'd1     , -6'd2     ,  6'd2     ,  6'd2     , -6'd1     , -6'd2     ,  6'd2     ,  6'd4     , -6'd2     , -6'd2     ,  6'd4     ,  6'd2     , -6'd2     , -6'd1      },
    '{  6'd0     ,  6'd6     , -6'd6     ,  6'd2     , -6'd6     ,  6'd2     ,  6'd2     ,  6'd4     , -6'd8     ,  6'd0     ,  6'd0     ,  6'd6     ,  6'd2     , -6'd6     ,  6'd2     ,  6'd0     , -6'd4     ,  6'd4     , -6'd2     ,  6'd0     ,  6'd4     , -6'd4     , -6'd4     ,  6'd0     ,  6'd4     , -6'd2     , -6'd8     ,  6'd6     , -6'd2     ,  6'd4     ,  6'd2     , -6'd8     ,  6'd4     ,  6'd12    , -6'd4     , -6'd2     ,  6'd8     , -6'd8     ,  6'd2     ,  6'd0     ,  6'd6     , -6'd8     , -6'd4     , -6'd6     , -6'd6     , -6'd2     ,  6'd0     , -6'd2     ,  6'd4     ,  6'd8      },
    '{  6'd0     , -6'd6     ,  6'd0     , -6'd8     , -6'd4     , -6'd6     , -6'd4     ,  6'd0     , -6'd6     , -6'd10    , -6'd12    , -6'd4     , -6'd8     ,  6'd0     ,  6'd6     , -6'd6     , -6'd2     , -6'd2     ,  6'd0     , -6'd6     ,  6'd6     ,  6'd2     ,  6'd0     , -6'd6     , -6'd8     , -6'd2     ,  6'd4     ,  6'd6     , -6'd2     ,  6'd6     ,  6'd10    ,  6'd0     , -6'd6     , -6'd8     ,  6'd4     , -6'd6     , -6'd6     ,  6'd6     ,  6'd0     , -6'd4     , -6'd6     ,  6'd4     , -6'd2     ,  6'd2     , -6'd2     ,  6'd4     ,  6'd0     , -6'd6     , -6'd6     , -6'd8      },
    '{  6'd0     , -6'd4     , -6'd4     ,  6'd0     ,  6'd4     ,  6'd2     , -6'd6     ,  6'd2     , -6'd2     ,  6'd2     ,  6'd2     , -6'd2     ,  6'd4     ,  6'd4     ,  6'd4     ,  6'd0     , -6'd2     ,  6'd0     ,  6'd6     , -6'd4     , -6'd2     , -6'd4     ,  6'd4     ,  6'd6     ,  6'd0     , -6'd6     ,  6'd0     ,  6'd2     ,  6'd2     ,  6'd2     ,  6'd0     , -6'd2     ,  6'd2     ,  6'd8     , -6'd2     , -6'd2     ,  6'd2     ,  6'd0     ,  6'd6     , -6'd2     , -6'd4     ,  6'd6     ,  6'd2     ,  6'd0     ,  6'd2     ,  6'd2     , -6'd2     ,  6'd2     ,  6'd2     ,  6'd0      },
    '{  6'd0     ,  6'd2     ,  6'd4     ,  6'd8     , -6'd4     , -6'd6     ,  6'd2     ,  6'd2     ,  6'd0     , -6'd2     , -6'd2     , -6'd6     ,  6'd0     , -6'd4     , -6'd2     ,  6'd2     , -6'd2     , -6'd2     , -6'd2     , -6'd2     ,  6'd2     ,  6'd0     ,  6'd0     , -6'd2     , -6'd2     , -6'd4     ,  6'd2     ,  6'd10    , -6'd4     ,  6'd6     , -6'd4     , -6'd2     ,  6'd0     ,  6'd0     , -6'd4     ,  6'd0     ,  6'd0     , -6'd4     , -6'd2     ,  6'd6     ,  6'd4     , -6'd4     , -6'd2     , -6'd2     , -6'd2     ,  6'd4     , -6'd4     , -6'd2     ,  6'd0     ,  6'd4      },
    '{  6'd0     ,  6'd4     , -6'd2     ,  6'd0     ,  6'd0     , -6'd4     ,  6'd4     , -6'd2     , -6'd2     , -6'd2     ,  6'd2     , -6'd4     , -6'd2     ,  6'd2     ,  6'd2     , -6'd2     , -6'd4     , -6'd2     , -6'd6     , -6'd2     , -6'd2     ,  6'd0     ,  6'd4     , -6'd6     , -6'd6     ,  6'd14    ,  6'd2     , -6'd4     , -6'd2     , -6'd4     ,  6'd2     , -6'd2     , -6'd2     , -6'd4     ,  6'd2     , -6'd2     ,  6'd2     , -6'd2     , -6'd4     , -6'd10    , -6'd2     ,  6'd0     ,  6'd4     ,  6'd0     ,  6'd0     ,  6'd2     ,  6'd0     ,  6'd0     , -6'd6     ,  6'd2      },
    '{  6'd0     ,  6'd0     , -6'd6     ,  6'd4     ,  6'd4     , -6'd2     , -6'd2     , -6'd2     , -6'd6     , -6'd6     , -6'd4     ,  6'd0     , -6'd4     ,  6'd0     , -6'd6     , -6'd6     , -6'd8     , -6'd12    ,  6'd0     ,  6'd0     , -6'd6     , -6'd8     ,  6'd0     , -6'd4     , -6'd4     ,  6'd4     , -6'd4     , -6'd2     , -6'd6     ,  6'd0     ,  6'd4     ,  6'd8     ,  6'd10    ,  6'd12    , -6'd4     , -6'd2     , -6'd2     ,  6'd0     ,  6'd6     ,  6'd6     ,  6'd6     ,  6'd6     ,  6'd0     , -6'd4     ,  6'd4     ,  6'd8     ,  6'd6     ,  6'd6     ,  6'd0     ,  6'd4      }
  };

  assign weights_n2 = '{
     4'd6,
     4'd3,
    -4'd3,
     4'd2,
     4'd6,
    -4'd5,
     4'd1,
     4'd3,
     4'd3,
    -4'd5,
     4'd2
  };
endmodule
